module csr import riscv_cpu_pkg::*;
#(
) (
  input  logic clk_i,
  input  logic rst_ni
);

endmodule : csr