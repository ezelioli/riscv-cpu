package riscv_cpu_pkg;

  /////////////////////////
  //    REGISTER FILE    //
  /////////////////////////
  parameter ADDR_WIDTH = 5;
  parameter DATA_WIDTH = 32;

  parameter CSR_WIDTH = 16;

endpackage : riscv_cpu_pkg